module top_module(input in, output out);
    assign in = out;
endmodule
