module (output zero);

    assign zero = 1'b0;
    // write nothing return 0

endmodule
